/*  Structure:
 *  Module States:
 *    Receive matrix length
 *    Matrix small - read
 *    Matrix large - read (portion)
 *    